
module ResetInverter(input RESET_IN, output RESET_OUT);
endmodule
