module BUFG ( output O, input  I);
    //buf B1 (O, I);
endmodule
