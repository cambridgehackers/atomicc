module mkZynqTop( input  CLK, input  RST_N,
  inout  [14 : 0] DDR_Addr, inout  [2 : 0] DDR_BankAddr,
  inout  DDR_CAS_n, inout  DDR_CKE, inout  DDR_CS_n, inout  DDR_Clk_n, inout  DDR_Clk_p,
  inout  [3 : 0] DDR_DM, inout  [31 : 0] DDR_DQ,
  inout  [3 : 0] DDR_DQS_n, inout  [3 : 0] DDR_DQS_p,
  inout  DDR_DRSTB, inout  DDR_ODT, inout  DDR_RAS_n,
  inout  FIXED_IO_ddr_vrn, inout  FIXED_IO_ddr_vrp, inout  DDR_WEB, inout  [53 : 0] MIO,
  inout  FIXED_IO_ps_clk, inout  FIXED_IO_ps_porb, inout  FIXED_IO_ps_srstb);

  wire ps7_clockGen_clkout0buffer_O;
  wire ps7_clockGen_pll_CLKFBOUT, ps7_clockGen_pll_CLKOUT0, ps7_clockGen_pll_CLKOUT0B;
  wire ps7_fclk_0_c_O, ps7_freset_0_r_O;
  wire [3 : 0] ps7_ps7_foo_FCLKCLK, ps7_ps7_foo_FCLKRESETN, maxigp0ARLEN, maxigp0AWLEN;

  wire ps7_b2c_0_IN1, ps7_b2c_0_IN2, ps7_b2c_3_IN1, ps7_b2c_3_IN2, ps7_b2c_0_OUT1, ps7_b2c_0_OUT2;
  assign ps7_b2c_0_IN1 = ps7_ps7_foo_FCLKCLK[0] ;
  assign ps7_b2c_0_IN2 = ps7_ps7_foo_FCLKRESETN[0] ;
  assign ps7_b2c_3_IN1 = ps7_ps7_foo_FCLKCLK[3] ;
  assign ps7_b2c_3_IN2 = ps7_ps7_foo_FCLKRESETN[3] ;
  CONNECTNET2 ps7_b2c_0(.IN1(ps7_b2c_0_IN1), .IN2(ps7_b2c_0_IN2), .OUT1(ps7_b2c_0_OUT1), .OUT2(ps7_b2c_0_OUT2));
  BUFG ps7_fclk_0_c(.I(ps7_b2c_0_OUT1), .O(ps7_fclk_0_c_O));
  BUFG ps7_freset_0_r(.I(ps7_b2c_0_OUT2), .O(ps7_freset_0_r_O));
  BUFG ps7_clockGen_clkout0buffer(.I(ps7_clockGen_pll_CLKOUT0), .O(ps7_clockGen_clkout0buffer_O));
  wire ps7_clockGen_pll_clkfbbuf_O, ps7_clockGen_pll_reset_RESET_OUT;
/* verilator lint_off PINMISSING */
  MMCME2_ADV #(.BANDWIDTH("OPTIMIZED"), .CLKFBOUT_USE_FINE_PS("FALSE"), .CLKOUT0_USE_FINE_PS("FALSE"),
        .CLKOUT1_USE_FINE_PS("FALSE"), .CLKOUT2_USE_FINE_PS("FALSE"), .CLKOUT3_USE_FINE_PS("FALSE"),
        .CLKOUT4_CASCADE("FALSE"), .CLKOUT4_USE_FINE_PS("FALSE"), .CLKOUT5_USE_FINE_PS("FALSE"),
        .CLKOUT6_USE_FINE_PS("FALSE"), .COMPENSATION("ZHOLD"), .STARTUP_WAIT("FALSE"),
        .CLKFBOUT_MULT_F(10.0), .CLKFBOUT_PHASE(0.0), .CLKIN1_PERIOD(10.0),
        .CLKIN2_PERIOD(0.0), .DIVCLK_DIVIDE(32'd1), .CLKOUT0_DIVIDE_F(5.0),
        .CLKOUT0_DUTY_CYCLE(0.5), .CLKOUT0_PHASE(0.0), .CLKOUT1_DIVIDE(32'd10),
        .CLKOUT1_DUTY_CYCLE(0.5), .CLKOUT1_PHASE(0.0), .CLKOUT2_DIVIDE(32'd10),
        .CLKOUT2_DUTY_CYCLE(0.5), .CLKOUT2_PHASE(0.0), .CLKOUT3_DIVIDE(32'd10),
        .CLKOUT3_DUTY_CYCLE(0.5), .CLKOUT3_PHASE(0.0), .CLKOUT4_DIVIDE(32'd10),
        .CLKOUT4_DUTY_CYCLE(0.5), .CLKOUT4_PHASE(0.0), .CLKOUT5_DIVIDE(32'd10),
        .CLKOUT5_DUTY_CYCLE(0.5), .CLKOUT5_PHASE(0.0), .CLKOUT6_DIVIDE(32'd10),
        .CLKOUT6_DUTY_CYCLE(0.5), .CLKOUT6_PHASE(0.0), .REF_JITTER1(1.0e-2),
        .REF_JITTER2(1.0e-2)) ps7_clockGen_pll(.CLKIN1(ps7_fclk_0_c_O),
        .RST(ps7_clockGen_pll_reset_RESET_OUT), .CLKIN2(1'd0), .CLKINSEL(1'd1),
        .DADDR(7'd0), .DCLK(1'd0), .DEN(1'd0), .DI(16'd0), .DWE(1'd0), .PSCLK(1'd0),
        .PSEN(1'd0), .PSINCDEC(1'd0), .PWRDWN(1'd0), .CLKFBIN(ps7_clockGen_pll_clkfbbuf_O), .LOCKED(),
        .CLKFBOUT(ps7_clockGen_pll_CLKFBOUT), .CLKFBOUTB(),
        .CLKOUT0(ps7_clockGen_pll_CLKOUT0), .CLKOUT0B(ps7_clockGen_pll_CLKOUT0B),
        .CLKOUT1(), .CLKOUT1B(), .CLKOUT2(), .CLKOUT2B(), .CLKOUT3(), .CLKOUT3B(),
        .CLKOUT4(), .CLKOUT5(), .CLKOUT6());
/* verilator lint_on PINMISSING */
  BUFG ps7_clockGen_pll_clkfbbuf(.I(ps7_clockGen_pll_CLKFBOUT), .O(ps7_clockGen_pll_clkfbbuf_O));
  ResetInverter ps7_clockGen_pll_reset(.RESET_IN(ps7_freset_0_r_O), .RESET_OUT(ps7_clockGen_pll_reset_RESET_OUT));

  wire [31 : 0] maxigp0ARADDR, maxigp0AWADDR, maxigp0WDATA;
  wire [11 : 0] maxigp0ARID, maxigp0AWID, maxigp0WID;
  wire maxigp0ARVALID, maxigp0AWVALID, maxigp0RREADY, maxigp0BREADY, maxigp0WLAST, maxigp0WVALID;
  wire maxigp0AWREADY, maxigp0WREADY, maxigp0BVALID, maxigp0ARREADY, maxigp0RVALID;
  wire [46 : 0] maxigp0RDATA;
  wire [13 : 0] maxigp0BRESP;
  wire ts_0_interrupt_0__read;
/* verilator lint_off PINMISSING */
  PS7 ps7_ps7_foo(.MAXIGP0ACLK(ps7_fclk_0_c_O),
        .MAXIGP1ACLK(ps7_fclk_0_c_O), .SAXIACPACLK(ps7_fclk_0_c_O), .SAXIGP0ACLK(ps7_fclk_0_c_O),
        .SAXIGP1ACLK(ps7_fclk_0_c_O), .SAXIHP0ACLK(ps7_fclk_0_c_O), .SAXIHP1ACLK(ps7_fclk_0_c_O),
        .SAXIHP2ACLK(ps7_fclk_0_c_O), .SAXIHP3ACLK(ps7_fclk_0_c_O),
        .DDRARB(0), .EMIOGPIOI(0), .EMIOI2C0SCLI(0), .EMIOI2C0SDAI(0), .EMIOI2C1SCLI(0),
        .EMIOI2C1SDAI(0), .EMIOSRAMINTIN(0), .EVENTEVENTI(0), .FCLKCLKTRIGN(0), .FPGAIDLEN(1),
        .IRQF2P({ 19'b0, ts_0_interrupt_0__read}),

        .MAXIGP0ARADDR(maxigp0ARADDR), .MAXIGP0ARID(maxigp0ARID), .MAXIGP0ARLEN(maxigp0ARLEN),
        .MAXIGP0ARVALID(maxigp0ARVALID), .MAXIGP0ARREADY(maxigp0ARREADY),

        .MAXIGP0RDATA(maxigp0RDATA[46:15]), .MAXIGP0RRESP(maxigp0RDATA[14:13]), .MAXIGP0RLAST(maxigp0RDATA[12]),
        .MAXIGP0RID(maxigp0RDATA[11:0]), .MAXIGP0RREADY(maxigp0RREADY), .MAXIGP0RVALID(maxigp0RVALID),

        .MAXIGP0AWADDR(maxigp0AWADDR), .MAXIGP0AWID(maxigp0AWID), .MAXIGP0AWLEN(maxigp0AWLEN),
        .MAXIGP0AWVALID(maxigp0AWVALID), .MAXIGP0AWREADY(maxigp0AWREADY),

        .MAXIGP0WDATA(maxigp0WDATA), .MAXIGP0WID(maxigp0WID), .MAXIGP0WLAST(maxigp0WLAST),
        .MAXIGP0WVALID(maxigp0WVALID), .MAXIGP0WREADY(maxigp0WREADY),

        .MAXIGP0BRESP(maxigp0BRESP[13:12]), .MAXIGP0BID(maxigp0BRESP[11:0]),
        .MAXIGP0BVALID(maxigp0BVALID), .MAXIGP0BREADY(maxigp0BREADY),
        .MAXIGP0ARBURST(), .MAXIGP0ARCACHE(), .MAXIGP0ARESETN(),
        .MAXIGP0ARLOCK(), .MAXIGP0ARPROT(), .MAXIGP0ARQOS(), .MAXIGP0ARSIZE(),
        .MAXIGP0AWBURST(), .MAXIGP0AWCACHE(), .MAXIGP0AWLOCK(), .MAXIGP0AWPROT(),
        .MAXIGP0AWQOS(), .MAXIGP0AWSIZE(), .MAXIGP0WSTRB(),

        .MAXIGP1ARREADY(0), .MAXIGP1AWREADY(0), .MAXIGP1BID(0), .MAXIGP1BRESP(0), .MAXIGP1BVALID(0),
        .MAXIGP1RDATA(0), .MAXIGP1RID(0), .MAXIGP1RLAST(0), .MAXIGP1RRESP(0), .MAXIGP1RVALID(0), .MAXIGP1WREADY(0),
        .SAXIACPARADDR(0), .SAXIACPARBURST(0), .SAXIACPARCACHE(0), .SAXIACPARID(0), .SAXIACPARLEN(0),
        .SAXIACPARLOCK(0), .SAXIACPARPROT(0), .SAXIACPARQOS(0), .SAXIACPARSIZE(0), .SAXIACPARUSER(0),
        .SAXIACPARVALID(0), .SAXIACPAWADDR(0), .SAXIACPAWBURST(0), .SAXIACPAWCACHE(0), .SAXIACPAWID(0),
        .SAXIACPAWLEN(0), .SAXIACPAWLOCK(0), .SAXIACPAWPROT(0), .SAXIACPAWQOS(0), .SAXIACPAWSIZE(0),
        .SAXIACPAWUSER(0), .SAXIACPAWVALID(0), .SAXIACPBREADY(0), .SAXIACPRREADY(0), .SAXIACPWDATA(0),
        .SAXIACPWID(0), .SAXIACPWLAST(0), .SAXIACPWSTRB(0), .SAXIACPWVALID(0),
        .SAXIGP0ARADDR(0), .SAXIGP0ARBURST(0), .SAXIGP0ARCACHE(0), .SAXIGP0ARID(0),
        .SAXIGP0ARLEN(0), .SAXIGP0ARLOCK(0), .SAXIGP0ARPROT(0), .SAXIGP0ARQOS(0),
        .SAXIGP0ARSIZE(0), .SAXIGP0ARVALID(0), .SAXIGP0AWADDR(0), .SAXIGP0AWBURST(0),
        .SAXIGP0AWCACHE(0), .SAXIGP0AWID(0), .SAXIGP0AWLEN(0), .SAXIGP0AWLOCK(0),
        .SAXIGP0AWPROT(0), .SAXIGP0AWQOS(0), .SAXIGP0AWSIZE(0), .SAXIGP0AWVALID(0),
        .SAXIGP0BREADY(0), .SAXIGP0RREADY(0), .SAXIGP0WDATA(0), .SAXIGP0WID(0),
        .SAXIGP0WLAST(0), .SAXIGP0WSTRB(0), .SAXIGP0WVALID(0), .SAXIGP1ARADDR(0),
        .SAXIGP1ARBURST(0), .SAXIGP1ARCACHE(0), .SAXIGP1ARID(0), .SAXIGP1ARLEN(0),
        .SAXIGP1ARLOCK(0), .SAXIGP1ARPROT(0), .SAXIGP1ARQOS(0), .SAXIGP1ARSIZE(0),
        .SAXIGP1ARVALID(0), .SAXIGP1AWADDR(0), .SAXIGP1AWBURST(0), .SAXIGP1AWCACHE(0),
        .SAXIGP1AWID(0), .SAXIGP1AWLEN(0), .SAXIGP1AWLOCK(0), .SAXIGP1AWPROT(0),
        .SAXIGP1AWQOS(0), .SAXIGP1AWSIZE(0), .SAXIGP1AWVALID(0), .SAXIGP1BREADY(0),
        .SAXIGP1RREADY(0), .SAXIGP1WDATA(0), .SAXIGP1WID(0), .SAXIGP1WLAST(0),
        .SAXIGP1WSTRB(0), .SAXIGP1WVALID(0), .SAXIHP0ARADDR(0), .SAXIHP0ARBURST(0),
        .SAXIHP0ARCACHE(0), .SAXIHP0ARID(0), .SAXIHP0ARLEN(0), .SAXIHP0ARLOCK(0),
        .SAXIHP0ARPROT(0), .SAXIHP0ARQOS(0), .SAXIHP0ARSIZE(0), .SAXIHP0ARVALID(0),
        .SAXIHP0AWADDR(0), .SAXIHP0AWBURST(0), .SAXIHP0AWCACHE(0), .SAXIHP0AWID(0),
        .SAXIHP0AWLEN(0), .SAXIHP0AWLOCK(0), .SAXIHP0AWPROT(0), .SAXIHP0AWQOS(0),
        .SAXIHP0AWSIZE(0), .SAXIHP0AWVALID(0), .SAXIHP0BREADY(0), .SAXIHP0RDISSUECAP1EN(0),
        .SAXIHP0RREADY(0), .SAXIHP0WDATA(0), .SAXIHP0WID(0), .SAXIHP0WLAST(0),
        .SAXIHP0WRISSUECAP1EN(0), .SAXIHP0WSTRB(0), .SAXIHP0WVALID(0), .SAXIHP1ARADDR(0),
        .SAXIHP1ARBURST(0), .SAXIHP1ARCACHE(0), .SAXIHP1ARID(0), .SAXIHP1ARLEN(0),
        .SAXIHP1ARLOCK(0), .SAXIHP1ARPROT(0), .SAXIHP1ARQOS(0), .SAXIHP1ARSIZE(0),
        .SAXIHP1ARVALID(0), .SAXIHP1AWADDR(0), .SAXIHP1AWBURST(0), .SAXIHP1AWCACHE(0),
        .SAXIHP1AWID(0), .SAXIHP1AWLEN(0), .SAXIHP1AWLOCK(0), .SAXIHP1AWPROT(0),
        .SAXIHP1AWQOS(0), .SAXIHP1AWSIZE(0), .SAXIHP1AWVALID(0), .SAXIHP1BREADY(0),
        .SAXIHP1RDISSUECAP1EN(0), .SAXIHP1RREADY(0), .SAXIHP1WDATA(0), .SAXIHP1WID(0),
        .SAXIHP1WLAST(0), .SAXIHP1WRISSUECAP1EN(0), .SAXIHP1WSTRB(0), .SAXIHP1WVALID(0),
        .SAXIHP2ARADDR(0), .SAXIHP2ARBURST(0), .SAXIHP2ARCACHE(0), .SAXIHP2ARID(0),
        .SAXIHP2ARLEN(0), .SAXIHP2ARLOCK(0), .SAXIHP2ARPROT(0), .SAXIHP2ARQOS(0),
        .SAXIHP2ARSIZE(0), .SAXIHP2ARVALID(0), .SAXIHP2AWADDR(0), .SAXIHP2AWBURST(0),
        .SAXIHP2AWCACHE(0), .SAXIHP2AWID(0), .SAXIHP2AWLEN(0), .SAXIHP2AWLOCK(0),
        .SAXIHP2AWPROT(0), .SAXIHP2AWQOS(0), .SAXIHP2AWSIZE(0), .SAXIHP2AWVALID(0),
        .SAXIHP2BREADY(0), .SAXIHP2RDISSUECAP1EN(0), .SAXIHP2RREADY(0), .SAXIHP2WDATA(0),
        .SAXIHP2WID(0), .SAXIHP2WLAST(0), .SAXIHP2WRISSUECAP1EN(0), .SAXIHP2WSTRB(0),
        .SAXIHP2WVALID(0), .SAXIHP3ARADDR(0), .SAXIHP3ARBURST(0), .SAXIHP3ARCACHE(0),
        .SAXIHP3ARID(0), .SAXIHP3ARLEN(0), .SAXIHP3ARLOCK(0), .SAXIHP3ARPROT(0),
        .SAXIHP3ARQOS(0), .SAXIHP3ARSIZE(0), .SAXIHP3ARVALID(0), .SAXIHP3AWADDR(0),
        .SAXIHP3AWBURST(0), .SAXIHP3AWCACHE(0), .SAXIHP3AWID(0), .SAXIHP3AWLEN(0),
        .SAXIHP3AWLOCK(0), .SAXIHP3AWPROT(0), .SAXIHP3AWQOS(0), .SAXIHP3AWSIZE(0),
        .SAXIHP3AWVALID(0), .SAXIHP3BREADY(0), .SAXIHP3RDISSUECAP1EN(0), .SAXIHP3RREADY(0),
        .SAXIHP3WDATA(0), .SAXIHP3WID(0), .SAXIHP3WLAST(0), .SAXIHP3WRISSUECAP1EN(0),
        .SAXIHP3WSTRB(0), .SAXIHP3WVALID(0), .EMIOGPIOO(), .EMIOGPIOTN(),
        .EMIOI2C0SCLO(), .EMIOI2C0SCLTN(), .EMIOI2C0SDAO(), .EMIOI2C0SDATN(),
        .EMIOI2C1SCLO(), .EMIOI2C1SCLTN(), .EMIOI2C1SDAO(), .EMIOI2C1SDATN(),
        .EVENTEVENTO(), .EVENTSTANDBYWFE(), .EVENTSTANDBYWFI(), .IRQP2F(),
        .MAXIGP1ARADDR(), .MAXIGP1ARBURST(), .MAXIGP1ARCACHE(), .MAXIGP1ARESETN(),
        .MAXIGP1ARID(), .MAXIGP1ARLEN(), .MAXIGP1ARLOCK(), .MAXIGP1ARPROT(),
        .MAXIGP1ARQOS(), .MAXIGP1ARSIZE(), .MAXIGP1ARVALID(), .MAXIGP1AWADDR(),
        .MAXIGP1AWBURST(), .MAXIGP1AWCACHE(), .MAXIGP1AWID(), .MAXIGP1AWLEN(),
        .MAXIGP1AWLOCK(), .MAXIGP1AWPROT(), .MAXIGP1AWQOS(), .MAXIGP1AWSIZE(),
        .MAXIGP1AWVALID(), .MAXIGP1BREADY(), .MAXIGP1RREADY(), .MAXIGP1WDATA(),
        .MAXIGP1WID(), .MAXIGP1WLAST(), .MAXIGP1WSTRB(), .MAXIGP1WVALID(),
        .SAXIACPARESETN(), .SAXIACPARREADY(), .SAXIACPAWREADY(), .SAXIACPBID(),
        .SAXIACPBRESP(), .SAXIACPBVALID(), .SAXIACPRDATA(), .SAXIACPRID(),
        .SAXIACPRLAST(), .SAXIACPRRESP(), .SAXIACPRVALID(), .SAXIACPWREADY(),
        .SAXIGP0ARESETN(), .SAXIGP0ARREADY(), .SAXIGP0AWREADY(), .SAXIGP0BID(),
        .SAXIGP0BRESP(), .SAXIGP0BVALID(), .SAXIGP0RDATA(), .SAXIGP0RID(),
        .SAXIGP0RLAST(), .SAXIGP0RRESP(), .SAXIGP0RVALID(), .SAXIGP0WREADY(),
        .SAXIGP1ARESETN(), .SAXIGP1ARREADY(), .SAXIGP1AWREADY(), .SAXIGP1BID(),
        .SAXIGP1BRESP(), .SAXIGP1BVALID(), .SAXIGP1RDATA(), .SAXIGP1RID(),
        .SAXIGP1RLAST(), .SAXIGP1RRESP(), .SAXIGP1RVALID(), .SAXIGP1WREADY(),
        .SAXIHP0ARESETN(), .SAXIHP0ARREADY(), .SAXIHP0AWREADY(), .SAXIHP0BID(),
        .SAXIHP0BRESP(), .SAXIHP0BVALID(), .SAXIHP0RDATA(), .SAXIHP0RID(),
        .SAXIHP0RLAST(), .SAXIHP0RRESP(), .SAXIHP0RVALID(), .SAXIHP0RACOUNT(),
        .SAXIHP0RCOUNT(), .SAXIHP0WACOUNT(), .SAXIHP0WCOUNT(), .SAXIHP0WREADY(),
        .SAXIHP1ARESETN(), .SAXIHP1ARREADY(), .SAXIHP1AWREADY(), .SAXIHP1BID(),
        .SAXIHP1BRESP(), .SAXIHP1BVALID(), .SAXIHP1RDATA(), .SAXIHP1RID(),
        .SAXIHP1RLAST(), .SAXIHP1RRESP(), .SAXIHP1RVALID(), .SAXIHP1RACOUNT(),
        .SAXIHP1RCOUNT(), .SAXIHP1WACOUNT(), .SAXIHP1WCOUNT(), .SAXIHP1WREADY(),
        .SAXIHP2ARESETN(), .SAXIHP2ARREADY(), .SAXIHP2AWREADY(), .SAXIHP2BID(),
        .SAXIHP2BRESP(), .SAXIHP2BVALID(), .SAXIHP2RDATA(), .SAXIHP2RID(),
        .SAXIHP2RLAST(), .SAXIHP2RRESP(), .SAXIHP2RVALID(), .SAXIHP2RACOUNT(),
        .SAXIHP2RCOUNT(), .SAXIHP2WACOUNT(), .SAXIHP2WCOUNT(), .SAXIHP2WREADY(),
        .SAXIHP3ARESETN(), .SAXIHP3ARREADY(), .SAXIHP3AWREADY(), .SAXIHP3BID(),
        .SAXIHP3BRESP(), .SAXIHP3BVALID(), .SAXIHP3RDATA(), .SAXIHP3RID(),
        .SAXIHP3RLAST(), .SAXIHP3RRESP(), .SAXIHP3RVALID(), .SAXIHP3RACOUNT(),
        .SAXIHP3RCOUNT(), .SAXIHP3WACOUNT(), .SAXIHP3WCOUNT(), .SAXIHP3WREADY(),
        .FCLKCLK(ps7_ps7_foo_FCLKCLK), .FCLKRESETN(ps7_ps7_foo_FCLKRESETN),
        .DDRA(DDR_Addr), .DDRBA(DDR_BankAddr), .DDRCASB(DDR_CAS_n),
        .DDRCKE(DDR_CKE), .DDRCKN(DDR_Clk_n), .DDRCKP(DDR_Clk_p),
        .DDRCSB(DDR_CS_n), .DDRDM(DDR_DM), .DDRDQ(DDR_DQ),
        .DDRDQSN(DDR_DQS_n), .DDRDQSP(DDR_DQS_p), .DDRDRSTB(DDR_DRSTB),
        .DDRODT(DDR_ODT), .DDRRASB(DDR_RAS_n), .DDRVRN(FIXED_IO_ddr_vrn),
        .DDRVRP(FIXED_IO_ddr_vrp), .DDRWEB(DDR_WEB), .PSCLK(FIXED_IO_ps_clk),
        .PSPORB(FIXED_IO_ps_porb), .PSSRSTB(FIXED_IO_ps_srstb), .MIO(MIO));
/* verilator lint_on PINMISSING */

  wire [38 : 0] ts_0_SRSData, ts_0_SWSData;
  wire [33 : 0] ts_0_SRSReq, ts_0_SWSReq;
  wire [5 : 0] ts_0_SWSDone;
  wire ts_0_RDY_SRSData, ts_0_RDY_SRSReq, ts_0_RDY_SWSData, ts_0_RDY_SWSDone, ts_0_RDY_SWSReq;
  wire RULE_SWSReq, RULEwriteDone, RULEwriteData;
  wire bufferAws_EMPTY_N, bufferAws_FULL_N, bufferWData_EMPTY_N, bufferWData_FULL_N, bufferBdone_FULL_N, readResp_FULL_N;
  assign RULEwriteDone = !maxigp0BVALID && ts_0_RDY_SWSDone ;
  assign RULE_SWSReq = bufferAws_EMPTY_N && ts_0_RDY_SWSReq ;
  assign RULEwriteData = bufferWData_EMPTY_N && ts_0_RDY_SWSData;
  assign maxigp0AWREADY = maxigp0AWVALID && !bufferAws_EMPTY_N;
  assign maxigp0WREADY = maxigp0WVALID && !bufferWData_EMPTY_N;

  FIFO2 #(.width(14), .guarded(1)) bufferBdone(.RST(ps7_freset_0_r_O), .CLK(ps7_fclk_0_c_O), .CLR(0),
        .D_IN( { 8'd0, ts_0_SWSDone }), .ENQ(RULEwriteDone),
        .D_OUT(maxigp0BRESP), .DEQ(maxigp0BVALID && maxigp0BREADY ),
        .FULL_N(bufferBdone_FULL_N), .EMPTY_N(maxigp0BVALID));
  FIFO1 #(.width(34), .guarded(1)) bufferAws(.RST(ps7_freset_0_r_O), .CLK(ps7_fclk_0_c_O), .CLR(0),
        .D_IN({ maxigp0AWADDR[17:0], { 4'd0, maxigp0AWLEN + 4'd1, 2'd0 }, maxigp0AWID[5:0] }), .ENQ(maxigp0AWREADY),
        .D_OUT(ts_0_SWSReq), .DEQ(RULE_SWSReq), .FULL_N(bufferAws_FULL_N), .EMPTY_N(bufferAws_EMPTY_N));
  FIFO2 #(.width(39), .guarded(1)) bufferWData(.RST(ps7_freset_0_r_O), .CLK(ps7_fclk_0_c_O), .CLR(0),
        .D_IN({maxigp0WDATA, maxigp0WID[5:0], maxigp0WLAST }), .ENQ(maxigp0WREADY),
        .D_OUT(ts_0_SWSData), .DEQ(RULEwriteData), .FULL_N(bufferWData_FULL_N), .EMPTY_N(bufferWData_EMPTY_N));

  wire bufferArs_EMPTY_N, bufferArs_FULL_N, RULE_SRSReq, RULE_getData;
  assign maxigp0ARREADY = maxigp0ARVALID && !bufferArs_EMPTY_N;
  assign RULE_SRSReq = bufferArs_EMPTY_N && ts_0_RDY_SRSReq ;
  assign RULE_getData = !maxigp0RVALID && ts_0_RDY_SRSData;

  FIFO1 #(.width(34), .guarded(1)) bufferArs(.RST(ps7_freset_0_r_O), .CLK(ps7_fclk_0_c_O), .CLR(0),
        .D_IN( { maxigp0ARADDR[17:0], { 4'd0, maxigp0ARLEN + 4'd1, 2'd0 }, maxigp0ARID[5:0] }), .ENQ(maxigp0ARREADY),
        .D_OUT(ts_0_SRSReq), .DEQ(RULE_SRSReq), .FULL_N(bufferArs_FULL_N), .EMPTY_N(bufferArs_EMPTY_N));
  FIFO2 #(.width(47), .guarded(1)) readResp(.RST(ps7_freset_0_r_O), .CLK(ps7_fclk_0_c_O), .CLR(0),
        .D_IN({ ts_0_SRSData[38:7], 9'd64, ts_0_SRSData[6:1] }), .ENQ(RULE_getData),
        .D_OUT(maxigp0RDATA), .DEQ(maxigp0RVALID && maxigp0RREADY), .FULL_N(readResp_FULL_N), .EMPTY_N(maxigp0RVALID));

  mkConnectalTop ts_0(.CLK(ps7_fclk_0_c_O), .RST_N(ps7_freset_0_r_O),
        .SRSReq(ts_0_SRSReq), .EN_SRSReq(RULE_SRSReq), .RDY_SRSReq(ts_0_RDY_SRSReq),
        .SRSData(ts_0_SRSData), .EN_SRSData(RULE_getData), .RDY_SRSData(ts_0_RDY_SRSData),
        .SWSReq(ts_0_SWSReq), .EN_SWSReq(RULE_SWSReq), .RDY_SWSReq(ts_0_RDY_SWSReq),
        .SWSData(ts_0_SWSData), .EN_SWSData(RULEwriteData), .RDY_SWSData(ts_0_RDY_SWSData),
        .SWSDone(ts_0_SWSDone), .EN_SWSDone(RULEwriteDone), .RDY_SWSDone(ts_0_RDY_SWSDone),
        .interrupt_0__read(ts_0_interrupt_0__read));
endmodule  // mkZynqTop
