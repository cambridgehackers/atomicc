../../../../atomicc-examples/examples/rulec/verilog/ProjectDefines.vh