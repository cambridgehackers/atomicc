../../../../atomicc-examples/examples/rulec/generated/rulec.generated.vh